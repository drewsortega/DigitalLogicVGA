module PS2_Input(
    input logic Clock,
    input logic Data,

    output logic Up,
    output logic Down,
    output logic Up,
    output logic Right
);

endmodule